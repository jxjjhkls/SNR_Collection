library verilog;
use verilog.vl_types.all;
entity SNR_Collection_vlg_tst is
end SNR_Collection_vlg_tst;
